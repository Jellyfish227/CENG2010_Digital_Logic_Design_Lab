library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
-- use IEEE.NUMERIC_STD.all;

entity ceng2010_hw1 is
    Port ( 
        clk : in STD_LOGIC;-- 100Mhz clk on Basys 3 FPGA board
        seg : out STD_LOGIC_VECTOR (6 downto 0);
        an : in STD_LOGIC_VECTOR (3 downto 0); -- 4 Anode signals
        dp : in std_logic := 1; --disabled decimal place
        btnC : in STD_LOGIC; --reset
        btnL : in STD_LOGIC; --rotate left
        btnR : in STD_LOGIC); --rotate right
end ceng2010_hw1;
the architecture Behavioral of ceng2010_hw1 is

signal displayed_number: STD_LOGIC_VECTOR (15 downto 0);
-- counting decimal number to be displayed on 4-digit 7-segment display
signal LED_BCD: STD_LOGIC_VECTOR (3 downto 0);
signal refresh_counter: STD_LOGIC_VECTOR (19 downto 0);
-- creating 10.5ms refresh period
signal LED_activating_counter: std_logic_vector(1 downto 0);
-- the other 2-bit for creating 4 LED-activating signals
-- count         0    ->  1  ->  2  ->  3
-- activates    LED1    LED2   LED3   LED4
-- and repeat
signal rst : std_logic;
signal first_digit : std_logic_vector(3 downto 0);
signal second_digit : std_logic_vector(3 downto 0);
signal third_digit : std_logic_vector(3 downto 0);
signal fourth_digit : std_logic_vector(3 downto 0);
signal state : std_logic_vector(1 downto 0):= "00";

begin 

    rst <= btnC;

    STATE_DETERMINE : process(btnC, btnL, btnR)
    begin
        if (rising_edge (btnR))
        
        end if;
    end process;
    
    -- VHDL code for BCD to 7-segment decoder
    -- Cathode patterns of the 7-segment LED display 
    process(LED_BCD)
    begin
        case LED_BCD is
        when "0000" => LED_out <= "0000001"; -- "0"     
        when "0001" => LED_out <= "1001111"; -- "1" 
        when "0010" => LED_out <= "0010010"; -- "2" 
        when "0011" => LED_out <= "0000110"; -- "3" 
        when "0100" => LED_out <= "1001100"; -- "4" 
        when "0101" => LED_out <= "0100100"; -- "5" 
        when "0110" => LED_out <= "0100000"; -- "6" 
        when "0111" => LED_out <= "0001111"; -- "7" 
        when "1000" => LED_out <= "0000000"; -- "8"     
        when "1001" => LED_out <= "0000100"; -- "9" 
        when "1010" => LED_out <= "0000010"; -- a
        when "1011" => LED_out <= "1100000"; -- b
        when "1100" => LED_out <= "0110001"; -- C
        when "1101" => LED_out <= "1000010"; -- d
        when "1110" => LED_out <= "0110000"; -- E
        when "1111" => LED_out <= "0111000"; -- F
        end case;
    end process;
    
    -- 7-segment display controller
    -- generate refresh period of 10.5ms
    process(clk,rst)
    begin 
        if(rst='1') then
            refresh_counter <= (others => '0');
        elsif(rising_edge(clk)) then
            refresh_counter <= refresh_counter + 1;
        end if;
    end process;

    LED_activating_counter <= refresh_counter(19 downto 18);
    -- 4-to-1 MUX to generate anode activating signals for 4 LEDs 
    process(LED_activating_counter)
    begin
        case LED_activating_counter is
        when "00" =>
            an <= "0111"; 
            -- activate LED1 and Deactivate LED2, LED3, LED4
            LED_BCD <= displayed_number(15 downto 12); 
            -- the first hex digit of the 16-bit number
        when "01" =>
            an <= "1011"; 
            -- activate LED2 and Deactivate LED1, LED3, LED4
            LED_BCD <= displayed_number(11 downto 8);
            -- the second hex digit of the 16-bit number
        when "10" =>
            an <= "1101"; 
            -- activate LED3 and Deactivate LED2, LED1, LED4
            LED_BCD <= displayed_number(7 downto 4);
            -- the third hex digit of the 16-bit number
        when "11" =>
            an <= "1110"; 
            -- activate LED4 and Deactivate LED2, LED3, LED1
            LED_BCD <= displayed_number(3 downto 0);
            -- the fourth hex digit of the 16-bit number    
        end case;
    end process;

    displayed_number <= "0111100010011010";
        
    
end Behavioral;